** Profile: "SCHEMATIC1-Response"  [ C:\Users\emanu\Desktop\DCE-GRUPO10\REALIMENTADOR\PSpice\Calculo-PSpiceFiles\SCHEMATIC1\Response.sim ] 

** Creating circuit file "Response.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of D:\Cadence\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.AC DEC 10000 1 10Meg
.OPTIONS ADVCONV
.OPTIONS SOLVER= 1
.OPTIONS METHOD= Default
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
